module signal_rename(
    input  sig_in,
    output sig_out
  );
  assign sig_out = sig_in;
endmodule
